-- megafunction wizard: %ALTSQRT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTSQRT 

-- ============================================================
-- File Name: altsqrt_varianceCalc.vhd
-- Megafunction Name(s):
-- 			ALTSQRT
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.1.0 Build 185 10/21/2015 SJ Lite Edition
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus Prime License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY altsqrt_varianceCalc IS
	PORT
	(
		clk		: IN STD_LOGIC ;
		radical		: IN STD_LOGIC_VECTOR (43 DOWNTO 0);
		q		: OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
		remainder		: OUT STD_LOGIC_VECTOR (22 DOWNTO 0)
	);
END altsqrt_varianceCalc;


ARCHITECTURE SYN OF altsqrt_variancecalc IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (21 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (22 DOWNTO 0);



	COMPONENT altsqrt
	GENERIC (
		pipeline		: NATURAL;
		q_port_width		: NATURAL;
		r_port_width		: NATURAL;
		width		: NATURAL;
		lpm_type		: STRING
	);
	PORT (
			clk	: IN STD_LOGIC ;
			radical	: IN STD_LOGIC_VECTOR (43 DOWNTO 0);
			q	: OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
			remainder	: OUT STD_LOGIC_VECTOR (22 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	q    <= sub_wire0(21 DOWNTO 0);
	remainder    <= sub_wire1(22 DOWNTO 0);

	ALTSQRT_component : ALTSQRT
	GENERIC MAP (
		pipeline => 11,
		q_port_width => 22,
		r_port_width => 23,
		width => 44,
		lpm_type => "ALTSQRT"
	)
	PORT MAP (
		clk => clk,
		radical => radical,
		q => sub_wire0,
		remainder => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "11"
-- Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "22"
-- Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "44"
-- Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL "clk"
-- Retrieval info: USED_PORT: q 0 0 22 0 OUTPUT NODEFVAL "q[21..0]"
-- Retrieval info: USED_PORT: radical 0 0 44 0 INPUT NODEFVAL "radical[43..0]"
-- Retrieval info: USED_PORT: remainder 0 0 23 0 OUTPUT NODEFVAL "remainder[22..0]"
-- Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
-- Retrieval info: CONNECT: @radical 0 0 44 0 radical 0 0 44 0
-- Retrieval info: CONNECT: q 0 0 22 0 @q 0 0 22 0
-- Retrieval info: CONNECT: remainder 0 0 23 0 @remainder 0 0 23 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_varianceCalc.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_varianceCalc.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_varianceCalc.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_varianceCalc.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altsqrt_varianceCalc_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
